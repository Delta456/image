module image
